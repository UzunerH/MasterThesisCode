`ifndef RV32_OPCODES
`define RV32_OPCODES

/*                            | func7 | rs2 | rs1 | 3 | rd  | op    | */
`define RV32_INSTR_LUI     32'b???????_?????_?????_???_?????_0110111 /* LUI */
`define RV32_INSTR_AUIPC   32'b???????_?????_?????_???_?????_0010111 /* AUIPC */
`define RV32_INSTR_JAL     32'b???????_?????_?????_???_?????_1101111 /* JAL */
`define RV32_INSTR_JALR    32'b???????_?????_?????_000_?????_1100111 /* JALR */
`define RV32_INSTR_BEQ     32'b???????_?????_?????_000_?????_1100011 /* BRANCH */
`define RV32_INSTR_BNE     32'b???????_?????_?????_001_?????_1100011
`define RV32_INSTR_BLT     32'b???????_?????_?????_100_?????_1100011
`define RV32_INSTR_BGE     32'b???????_?????_?????_101_?????_1100011
`define RV32_INSTR_BLTU    32'b???????_?????_?????_110_?????_1100011
`define RV32_INSTR_BGEU    32'b???????_?????_?????_111_?????_1100011
`define RV32_INSTR_LB      32'b???????_?????_?????_000_?????_0000011 /* LOAD */
`define RV32_INSTR_LH      32'b???????_?????_?????_001_?????_0000011
`define RV32_INSTR_LW      32'b???????_?????_?????_010_?????_0000011
`define RV32_INSTR_LBU     32'b???????_?????_?????_100_?????_0000011
`define RV32_INSTR_LHU     32'b???????_?????_?????_101_?????_0000011
`define RV32_INSTR_SB      32'b???????_?????_?????_000_?????_0100011 /* STORE */
`define RV32_INSTR_SH      32'b???????_?????_?????_001_?????_0100011
`define RV32_INSTR_SW      32'b???????_?????_?????_010_?????_0100011
`define RV32_INSTR_ADDI    32'b???????_?????_?????_000_?????_0010011 /* OP-IMM */
`define RV32_INSTR_SLTI    32'b???????_?????_?????_010_?????_0010011
`define RV32_INSTR_SLTIU   32'b???????_?????_?????_011_?????_0010011
`define RV32_INSTR_XORI    32'b???????_?????_?????_100_?????_0010011
`define RV32_INSTR_ORI     32'b???????_?????_?????_110_?????_0010011
`define RV32_INSTR_ANDI    32'b???????_?????_?????_111_?????_0010011
`define RV32_INSTR_SLLI    32'b0000000_?????_?????_001_?????_0010011
`define RV32_INSTR_SRLI    32'b0000000_?????_?????_101_?????_0010011
`define RV32_INSTR_SRAI    32'b0100000_?????_?????_101_?????_0010011
`define RV32_INSTR_ADD     32'b0000000_?????_?????_000_?????_0110011 /* OP */
`define RV32_INSTR_SUB     32'b0100000_?????_?????_000_?????_0110011
`define RV32_INSTR_SLL     32'b0000000_?????_?????_001_?????_0110011
`define RV32_INSTR_SLT     32'b0000000_?????_?????_010_?????_0110011
`define RV32_INSTR_SLTU    32'b0000000_?????_?????_011_?????_0110011
`define RV32_INSTR_XOR     32'b0000000_?????_?????_100_?????_0110011
`define RV32_INSTR_SRL     32'b0000000_?????_?????_101_?????_0110011
`define RV32_INSTR_SRA     32'b0100000_?????_?????_101_?????_0110011
`define RV32_INSTR_OR      32'b0000000_?????_?????_110_?????_0110011
`define RV32_INSTR_AND     32'b0000000_?????_?????_111_?????_0110011
`define RV32_INSTR_FENCE   32'b???????_?????_?????_000_?????_0001111 /* MISC-MEM */
`define RV32_INSTR_FENCE_I 32'b???????_?????_?????_001_?????_0001111
`define RV32_INSTR_ECALL   32'b0000000_00000_00000_000_00000_1110011 /* SYSTEM */
`define RV32_INSTR_EBREAK  32'b0000000_00001_00000_000_00000_1110011
`define RV32_INSTR_MRET    32'b0011000_00010_00000_000_00000_1110011
`define RV32_INSTR_WFI     32'b0001000_00101_00000_000_00000_1110011
`define RV32_INSTR_CSRRW   32'b???????_?????_?????_001_?????_1110011
`define RV32_INSTR_CSRRS   32'b???????_?????_?????_010_?????_1110011
`define RV32_INSTR_CSRRC   32'b???????_?????_?????_011_?????_1110011
`define RV32_INSTR_CSRRWI  32'b???????_?????_?????_101_?????_1110011
`define RV32_INSTR_CSRRSI   32'b???????_?????_?????_110_?????_1110011
`define RV32_INSTR_CSRRCI   32'b???????_?????_?????_111_?????_1110011
`define RV32_INSTR_NLD_NL    	32'b???????_?????_?????_???_?????_0000111 /* NLU-LOAD */
`define RV32_INSTR_NLD_L     	32'b???????_?????_?????_???_?????_0001011 
`define RV32_INSTR_NNL_ANF   	32'b0000000_00000_?????_000_?????_0011011 /* NLU-OPs */
`define RV32_INSTR_NNL_AES_E   	32'b0000000_00000_?????_001_?????_0011011 
`define RV32_INSTR_NNL_AES_D   	32'b0000000_00000_?????_010_?????_0011011 
`define RV32_INSTR_NMU 		 	32'b0000000_00000_?????_011_?????_0011011 
`define RV32_INSTR_NMA0 		32'b0000000_00000_?????_100_?????_0011011 
`define RV32_INSTR_NMA1 		32'b0000000_00000_?????_101_?????_0011011 
`define RV32_INSTR_NMA2 		32'b0000000_00000_?????_110_?????_0011011 
`define RV32_INSTR_NMA3 		32'b0000000_00000_?????_111_?????_0011011 


`define RV32_INSTR_NOP     32'b0000000_00000_00000_000_00000_0010011

`define RV32_OPCODE_JAL    7'b1101111
`define RV32_OPCODE_BRANCH 7'b1100011

`endif
